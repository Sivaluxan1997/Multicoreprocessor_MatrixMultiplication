module ins_memory(clk,addr1,addr2,addr3,addr4,ins_out1,ins_out2,ins_out3,ins_out4,im_write_en,im_input_data,im_addr);
//module im(clk,write_en,addr,ins_in,ins_out);
	input clk;
	//input write_en;  //we can remove write_en and ins_in
	input [15:0] addr1,addr2,addr3,addr4;
	//input [15:0] ins_in;
	output reg [15:0] ins_out1,ins_out2,ins_out3,ins_out4;
	input im_write_en;
   input [15:0] im_input_data;
   input [15:0] im_addr;
	
	reg [15:0] ins_ram[100:0];
	
	/*parameter
	clall= 16'd3,
	nop=16'd4,
	ldac=16'd5,
	mvacti=16'd7,
	mvactj=16'd8,
	mvactk=16'd9,
	mvactr=16'd10,
	mvactar=16'd11,
	mvacr=16'd12,
	mvacao=16'd13,
	mvacdar=16'd14,
	mvace=16'd15,
	mvtiac=16'd16,
	mvtjac=16'd17,
	mvtkac=16'd18,
	mvrac=16'd19,
	add=16'd20,
	mul=16'd21,
	sub=16'd22,
	incac=16'd23,
	incri=16'd24,
	incrj=16'd25,
	incrk=16'd26,
	incao=16'd27,
	stac=16'd28,
	jumpnz=16'd29,
	mvtarr=16'd33,
	mver=16'd34,
	mvtrr=16'd35,
	mvrir=16'd36,
	mvrjr=16'd37,
	mvrkr=16'd38,
	clac=16'd39,
	clri=16'd40,
	clrj=16'd41,
	clrk=16'd42,
	mvaodar=16'd43,
	core_en=16'd49,
	mvaor=16'd50,
	jumpz=16'd51,
	endop=16'd44;*/
	
	initial begin
	//4 core
		/*ram[0]=clall;
		ram[1]=ldac;
		ram[2]=mvacti;
		ram[3]=ldac;
		ram[4]=mvactj;
		ram[5]=ldac;
		ram[6]=mvactk;
		ram[7]=core_en;
		ram[8]=core_en;
		ram[9]=core_en;
		ram[10]=mvtiac;
		ram[11]=mvacr;
		ram[12]=mvtjac;
		ram[13]=mul;
		ram[14]=mvactar;
		ram[15]=mvtjac;
		ram[16]=mvacr;
		ram[17]=mvtkac;
		ram[18]=mul;
		ram[19]=mvtarr;
		ram[20]=add;
		ram[21]=incac;
		ram[22]=incac;
		ram[23]=incac;
		ram[24]=mvacao;
		ram[25]=mvrir;  //loop2.....loop1.....loop3
		ram[26]=mvtjac;
		ram[27]=mul;
		ram[28]=mvrjr;
		ram[29]=add;
		ram[30]=incac;
		ram[31]=incac;
		ram[32]=incac;
		ram[33]=mvacdar;
		ram[34]=ldac;
		ram[35]=mvace;
		ram[36]=mvtkac;
		ram[37]=mul;
		ram[38]=mvrkr;
		ram[39]=add;
		ram[40]=mvtarr;
		ram[41]=add;
		ram[42]=incac;
		ram[43]=incac;
		ram[44]=incac;
		ram[45]=mvacdar;
		ram[46]=ldac;
		ram[47]=mver;
		ram[48]=mul;
		ram[49]=mvtrr;
		ram[50]=add;
		ram[51]=mvactr;
		ram[52]=incrj;
		ram[53]=mvrjr;
		ram[54]=mvtjac;
		ram[55]=sub;
		ram[56]=jumpnz;
		ram[57]=16'd25;//jump to loop2
		ram[58]=mvrir;
		ram[59]=mvtkac;
		ram[60]=mul;
		ram[61]=mvrkr;
		ram[62]=add;
		ram[63]=mvaor;
		ram[64]=add;
		ram[65]=mvacdar;
		ram[66]=mvtrr;
		ram[67]=mvrac;
		//ram[66]=mvaodar;
		ram[68]=stac;
		//ram[68]=incao;
		ram[69]=clac;
		ram[70]=mvactr;
		ram[71]=clrj;
		ram[72]=incrk;
		ram[73]=mvrkr;
		ram[74]=mvtkac;
		ram[75]=sub;
		ram[76]=jumpnz;
		ram[77]=16'd25;//jump to loop1
		ram[78]=clac;
		ram[79]=mvactr;
		ram[80]=clrj;
		ram[81]=clrk;
		ram[82]=incri;
		ram[83]=incri;
		ram[84]=incri;
		ram[85]=incri;
		ram[86]=mvrir;
		ram[87]=mvtiac;
		ram[88]=sub;
		ram[89]=jumpnz;
		ram[90]=16'd25;//jump to loop3
		ram[91]=endop;*/
		//3 core
		/*ram[0]=clall;
		ram[1]=ldac;
		ram[2]=mvacti;
		ram[3]=ldac;
		ram[4]=mvactj;
		ram[5]=ldac;
		ram[6]=mvactk;
		//ram[7]=core_en;
		ram[7]=core_en;
		ram[8]=core_en;
		ram[9]=mvtiac;
		ram[10]=mvacr;
		ram[11]=mvtjac;
		ram[12]=mul;
		ram[13]=mvactar;
		ram[14]=mvtjac;
		ram[15]=mvacr;
		ram[16]=mvtkac;
		ram[17]=mul;
		ram[18]=mvtarr;
		ram[19]=add;
		ram[20]=incac;
		ram[21]=incac;
		ram[22]=incac;
		ram[23]=mvacao;
		ram[24]=mvrir;  //loop2.....loop1.....loop3
		ram[25]=mvtjac;
		ram[26]=mul;
		ram[27]=mvrjr;
		ram[28]=add;
		ram[29]=incac;
		ram[30]=incac;
		ram[31]=incac;
		ram[32]=mvacdar;
		ram[33]=ldac;
		ram[34]=mvace;
		ram[35]=mvtkac;
		ram[36]=mul;
		ram[37]=mvrkr;
		ram[38]=add;
		ram[39]=mvtarr;
		ram[40]=add;
		ram[41]=incac;
		ram[42]=incac;
		ram[43]=incac;
		ram[44]=mvacdar;
		ram[45]=ldac;
		ram[46]=mver;
		ram[47]=mul;
		ram[48]=mvtrr;
		ram[49]=add;
		ram[50]=mvactr;
		ram[51]=incrj;
		ram[52]=mvrjr;
		ram[53]=mvtjac;
		ram[54]=sub;
		ram[55]=jumpnz;
		ram[56]=16'd24;//jump to loop2
		ram[57]=mvrir;
		ram[58]=mvtkac;
		ram[59]=mul;
		ram[60]=mvrkr;
		ram[61]=add;
		ram[62]=mvaor;
		ram[63]=add;
		ram[64]=mvacdar;
		ram[65]=mvtrr;
		ram[66]=mvrac;
		//ram[66]=mvaodar;
		ram[67]=stac;
		//ram[68]=incao;
		ram[68]=clac;
		ram[69]=mvactr;
		ram[70]=clrj;
		ram[71]=incrk;
		ram[72]=mvrkr;
		ram[73]=mvtkac;
		ram[74]=sub;
		ram[75]=jumpnz;
		ram[76]=16'd24;//jump to loop1
		ram[77]=clac;
		ram[78]=mvactr;
		ram[79]=clrj;
		ram[80]=clrk;
		ram[81]=incri;
		ram[82]=incri;
		ram[83]=incri;
		//ram[85]=incri;
		ram[84]=mvrir;
		ram[85]=mvtiac;
		ram[86]=sub;
		ram[87]=jumpnz;
		ram[88]=16'd24;//jump to loop3
		ram[89]=endop;*/
		//two core
		/*ram[0]=clall;
		ram[1]=ldac;
		ram[2]=mvacti;
		ram[3]=ldac;
		ram[4]=mvactj;
		ram[5]=ldac;
		ram[6]=mvactk;
		ram[7]=core_en;
		//ram[8]=incri;
		ram[8]=mvtiac;
		ram[9]=mvacr;
		ram[10]=mvtjac;
		ram[11]=mul;
		ram[12]=mvactar;
		ram[13]=mvtjac;
		ram[14]=mvacr;
		ram[15]=mvtkac;
		ram[16]=mul;
		ram[17]=mvtarr;
		ram[18]=add;
		ram[19]=incac;
		ram[20]=incac;
		ram[21]=incac;
		ram[22]=mvacao;
		ram[23]=mvrir;  //loop2.....loop1.....loop3
		ram[24]=mvtjac;
		ram[25]=mul;
		ram[26]=mvrjr;
		ram[27]=add;
		ram[28]=incac;
		ram[29]=incac;
		ram[30]=incac;
		ram[31]=mvacdar;
		ram[32]=ldac;
		ram[33]=mvace;
		ram[34]=mvtkac;
		ram[35]=mul;
		ram[36]=mvrkr;
		ram[37]=add;
		ram[38]=mvtarr;
		ram[39]=add;
		ram[40]=incac;
		ram[41]=incac;
		ram[42]=incac;
		ram[43]=mvacdar;
		ram[44]=ldac;
		ram[45]=mver;
		ram[46]=mul;
		ram[47]=mvtrr;
		ram[48]=add;
		ram[49]=mvactr;
		ram[50]=incrj;
		ram[51]=mvrjr;
		ram[52]=mvtjac;
		ram[53]=sub;
		ram[54]=jumpnz;
		ram[55]=16'd23;//jump to loop2
		ram[56]=mvrir;
		ram[57]=mvtkac;
		ram[58]=mul;
		ram[59]=mvrkr;
		ram[60]=add;
		ram[61]=mvaor;
		ram[62]=add;
		ram[63]=mvacdar;
		ram[64]=mvtrr;
		ram[65]=mvrac;
		//ram[66]=mvaodar;
		ram[66]=stac;
		//ram[68]=incao;
		ram[67]=clac;
		ram[68]=mvactr;
		ram[69]=clrj;
		ram[70]=incrk;
		ram[71]=mvrkr;
		ram[72]=mvtkac;
		ram[73]=sub;
		ram[74]=jumpnz;
		ram[75]=16'd23;//jump to loop1
		ram[76]=clac;
		ram[77]=mvactr;
		ram[78]=clrj;
		ram[79]=clrk;
		ram[80]=incri;
		ram[81]=incri;
		ram[82]=mvrir;
		ram[83]=mvtiac;
		ram[84]=sub;
		ram[85]=jumpnz;
		ram[86]=16'd23;//jump to loop3
		ram[87]=endop;*/
		//single core
		/*ram[0]=clall;
		ram[1]=ldac;
		ram[2]=mvacti;
		ram[3]=ldac;
		ram[4]=mvactj;
		ram[5]=ldac;
		ram[6]=mvactk;
		ram[7]=mvtiac;
		ram[8]=mvacr;
		ram[9]=mvtjac;
		ram[10]=mul;
		ram[11]=mvactar;
		ram[12]=mvtjac;
		ram[13]=mvacr;
		ram[14]=mvtkac;
		ram[15]=mul;
		ram[16]=mvtarr;
		ram[17]=add;
		ram[18]=incac;
		ram[19]=incac;
		ram[20]=incac;
		ram[21]=mvacao;
		ram[22]=mvrir;  //loop2.....loop1.....loop3
		ram[23]=mvtjac;
		ram[24]=mul;
		ram[25]=mvrjr;
		ram[26]=add;
		ram[27]=incac;
		ram[28]=incac;
		ram[29]=incac;
		ram[30]=mvacdar;
		ram[31]=ldac;
		ram[32]=mvace;
		ram[33]=mvtkac;
		ram[34]=mul;
		ram[35]=mvrkr;
		ram[36]=add;
		ram[37]=mvtarr;
		ram[38]=add;
		ram[39]=incac;
		ram[40]=incac;
		ram[41]=incac;
		ram[42]=mvacdar;
		ram[43]=ldac;
		ram[44]=mver;
		ram[45]=mul;
		ram[46]=mvtrr;
		ram[47]=add;
		ram[48]=mvactr;
		ram[49]=incrj;
		ram[50]=mvrjr;
		ram[51]=mvtjac;
		ram[52]=sub;
		ram[53]=jumpnz;
		ram[54]=16'd22;//jump to loop2
		ram[55]=mvtrr;
		ram[56]=mvrac;
		ram[57]=mvaodar;
		ram[58]=stac;
		ram[59]=incao;
		ram[60]=clac;
		ram[61]=mvactr;
		ram[62]=clrj;
		ram[63]=incrk;
		ram[64]=mvrkr;
		ram[65]=mvtkac;
		ram[66]=sub;
		ram[67]=jumpnz;
		ram[68]=16'd22;//jump to loop1
		ram[69]=clac;
		ram[70]=mvactr;
		ram[71]=clrj;
		ram[72]=clrk;
		ram[73]=incri;
		ram[74]=mvrir;
		ram[75]=mvtiac;
		ram[76]=sub;
		ram[77]=jumpnz;
		ram[78]=16'd22;//jump to loop3
		ram[79]=endop;*/
	end
	
	always @(posedge clk)
		begin
			//if (write_en==1)
				//ram[addr] <= ins_in[15:0];
			//else
			//if (addr1==addr2)
				ins_out1 <= ins_ram[addr1];
				ins_out2 <= ins_ram[addr2];
				ins_out3 <= ins_ram[addr3];
				ins_out4 <= ins_ram[addr4];
				
			if (im_write_en == 1) begin
				ins_ram[im_addr]<=im_input_data;
			end
					
			
		end
endmodule

	